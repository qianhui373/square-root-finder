




`timescale 1 ns/1 ns

module tb_newton();

 
endmodule